`define N = 4